
module system (
	clk_clk,
	sine_wave_generator_0_conduit_end_export,
	reset_reset_n);	

	input		clk_clk;
	output	[9:0]	sine_wave_generator_0_conduit_end_export;
	input		reset_reset_n;
endmodule
