
module system (
	clk_clk,
	reset_reset_n,
	sine_wave_generator_0_conduit_end_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[9:0]	sine_wave_generator_0_conduit_end_export;
endmodule
